module hello_world();
initial
$display("hello verilog world!");
endmodule
