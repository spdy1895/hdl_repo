`define TRUE 1'b1
`define FLASE 1'b0
`define Y2R_DELAY 3
`define R2G_ DELAY 2

module sig_control (
    
);

endmodule //sig_control
