module hello_world():
$display("hello verilog world!");
endmodule
